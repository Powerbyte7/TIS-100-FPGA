library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

entity tis_node_tb is
end entity;

architecture rtl of tis_node_tb is
    
begin
    t0 : work.tis_node port map ()
end architecture;